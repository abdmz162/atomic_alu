module memory()

endmodule